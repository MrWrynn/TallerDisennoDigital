module shift1bit (
		input logic In,
		output logic Out);
		
assign Out = In;
		
		
endmodule