module divisor #(N=4) (
				input logic [N-1:0] aIn,
				input logic [N-1:0] bIn,
				output logic [N-1:0] cOut,
				output logic [N-1:0] mod);



				
endmodule